********************************************************************************
* Library Name: Pipeline_ADC
* Cell Name: bootstrap
* View Name: schematic
********************************************************************************

.SUBCKT bootstrap vdd gnd vin out clk
XI0 clk clkb gnd vdd / inv_dac
MN1 n3 clkb gnd gnd n18 W=20u L=200n m=1
MP2 n2 n4 vdd vdd p18 W=20u L=200n m=1
MP4 n1 clk vdd vdd p18 W=20u L=200n m=1
MN4 n1 clk n3 gnd n18 W=20u L=200n m=1
MP1 n4 n1 n2 vdd p18 W=20u L=200n m=1
MN3 n1 n4 n3 gnd n18 W=20u L=200n m=1
MN5 n4 vdd n5 gnd n18 W=20u L=200n m=1
MN7 vin n4 n3 gnd n18 W=20u L=200n m=1
MP3 vin clkb n3 vdd p18 W=20u L=200n m=1
MP5 vdd clkb n5 vdd p18 W=20u L=200n m=1
MN6 n5 clkb gnd gnd n18 W=20u L=200n m=1
MNS out n4 vin gnd n18 W=20u L=200n m=1

Cb n2 n3 200f

.ENDS